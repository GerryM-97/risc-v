library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use WORK.generics.all;

ENTITY op_decoder IS
PORT ( 
		--input
		INSTRUCTION_IN 	: in instruction;
		
		--output
		INSTRUCTION_F 	: out instruction_format;
		OP_DECODED 		: out operation
);
END ENTITY;

ARCHITECTURE behav OF op_decoder IS

SIGNAL OP_DEC : operation;

BEGIN

OP_DECODED <= OP_DEC;

OP_DEC <=   	ADD 	WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0110011" AND INSTRUCTION_IN(14 DOWNTO 12) = "000" 	ELSE 	
				ADDI	WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0010011" AND INSTRUCTION_IN(14 DOWNTO 12) = "000"	ELSE
				AUIPC	WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0010111" 											ELSE
				LUI		WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0110111" 											ELSE
				BEQ		WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "1100011" AND INSTRUCTION_IN(14 DOWNTO 12) = "000"	ELSE
				LW		WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0000011" AND INSTRUCTION_IN(14 DOWNTO 12) = "010"	ELSE
				SRAI	WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0010011" AND INSTRUCTION_IN(14 DOWNTO 12) = "101"	ELSE
				ANDI	WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0010011" AND INSTRUCTION_IN(14 DOWNTO 12) = "111"	ELSE
				XOR_T	WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0110011" AND INSTRUCTION_IN(14 DOWNTO 12) = "100"	ELSE
				SLT		WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0110011" AND INSTRUCTION_IN(14 DOWNTO 12) = "010"	ELSE
				JAL		WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "1101111" 											ELSE
				SW		WHEN 		INSTRUCTION_IN(opcode_len-1 DOWNTO 0) = "0100011" AND INSTRUCTION_IN(14 DOWNTO 12) = "010"	ELSE
				ADDI; --NOP

instruction_f <= R_type 	WHEN OP_DEC = ADD OR OP_DEC = XOR_T ELSE
				 I_type 	WHEN OP_DEC = ADDI OR OP_DEC = LW OR OP_DEC = SRAI OR OP_DEC = ANDI OR OP_DEC = NOP ELSE
				 B_type 	WHEN OP_DEC = BEQ 	ELSE
				 S_type 	WHEN OP_DEC = SW ELSE
				 J_type 	WHEN OP_DEC = JAL ELSE
				 U_type 	WHEN OP_DEC = AUIPC OR OP_DEC = LUI ELSE
				 I_type; --nop operation

END ARCHITECTURE;
